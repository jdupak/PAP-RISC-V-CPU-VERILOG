module InstructionMemory(
    input wire[0:0] clk,
    input wire[31:0] read_idx,
    output reg[31:0] read_data
);
    reg[31:0] mem[128:0];

    always @ (read_idx) begin
        read_data = mem[read_idx[9:2]];
    end

    initial begin
        //read_data = 32'b000000000000_00000_000_00000_0010011; // NOP
        mem[0] = 32'b0000000_00000_00000_000_00000_0010011; // NOP
        mem[1] = 32'b0000010_00010_00001_001_01000_1100011;
        mem[2] = 32'b0000000_00010_00001_000_00001_0010011;
        mem[3] = 32'b0000000_00111_00001_000_00001_0010011;
        mem[4] = 32'b0000000_00001_00000_000_00000_0100011;
        mem[5] = 32'b0000000_00001_00001_000_00001_0010011;
        mem[6] = 32'b0000000_00011_00001_000_00001_0010011;
        mem[7] = 32'b0000000_00000_00000_000_00001_0000011;
        mem[8] = 32'b0000000_00101_00001_000_00010_0010011;
        mem[9] = 32'b1111111_00001_11111_111_00000_1101111;
        mem[10] =32'b0000000_00001_00000_000_00000_1110011; // BREAK
    end
endmodule
