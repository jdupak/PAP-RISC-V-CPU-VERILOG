module InstructionMemory(
    input wire[0:0] clk,
    input wire[31:0] read_idx,
    output reg[31:0] read_data
);
    reg[31:0] mem[128:0];
    integer fd, i;

    always @ (read_idx) begin
        read_data = mem[read_idx[9:2]];
    end

    initial begin
        fd = $fopen("gcd.bin","rb");
        i = $fread(mem, fd);
        $fclose(fd);
        // TEST
        //mem[0] = 32'b0000000_00000_00000_000_00000_0010011; // NOP
        //mem[1] = 32'b0000010_00010_00001_001_01000_1100011;
        //mem[2] = 32'b0000000_00010_00001_000_00001_0010011;
        //mem[3] = 32'b0000000_00111_00001_000_00001_0010011;
        //mem[4] = 32'b0000000_00001_00000_000_00000_0100011;
        //mem[5] = 32'b0000000_00001_00001_000_00001_0010011;
        //mem[6] = 32'b0000000_00011_00001_000_00001_0010011;
        //mem[7] = 32'b0000000_00000_00000_000_00001_0000011;
        //mem[8] = 32'b0000000_00101_00001_000_00010_0010011;
        //mem[9] = 32'b1111111_00001_11111_111_00000_1101111;
        //mem[10] =32'b0000000_00001_00000_000_00000_1110011; // BREAK

        // GCD
        //mem[0] = 32'b0000000_00000_00000_000_00000_0010011; // NOP
        //mem[1] = 32'b0000000_00100_00000_010_00001_0000011;
        //mem[2] = 32'b0000000_01000_00000_010_00010_0000011;
        //mem[3] = 32'b0000011_00001_00000_000_01000_1100011;
        //mem[4] = 32'b0000011_00010_00000_000_10000_1100011;
        //mem[5] = 32'b0000000_00000_00000_100_00100_0110011;
        //mem[6] = 32'b0000000_00010_00001_110_00011_0110011;
        //mem[7] = 32'b0000000_00001_00011_111_00011_0010011;
        //mem[8] = 32'b0000000_10000_00011_001_10100_1100011;
        //mem[9] = 32'b0000000_00001_00100_111_00100_0010011;
        //mem[10] = 32'b0000000_00001_00001_101_00001_0010011;
        //mem[11] = 32'b0000000_00001_00010_101_00010_0010011;
        //mem[12] = 32'b1111111_10101_11111_111_00000_1101111;
        //mem[13] = 32'b0000000_00001_00001_111_00011_0010011;
        //mem[14] = 32'b0000000_00011_00000_001_11000_1100011;
        //mem[15] = 32'b0000000_00001_00001_101_00001_0010011;
        //mem[16] = 32'b1111111_10101_11111_111_00000_1101111;
        //mem[17] = 32'b0000000_00001_00010_111_00011_0010011;
        //mem[18] = 32'b0000000_00011_00000_001_11000_1100011;
        //mem[19] = 32'b0000000_00001_00010_101_00010_0010011;
        //mem[20] = 32'b1111111_10101_11111_111_00000_1101111;
        //mem[21] = 32'b0000000_00000_00000_000_00000_0010011; // NOP
        //mem[22] = 32'b0000001_00011_00000_001_00000_1100011; //
        //mem[23] = 32'b0000000_00000_00001_100_00011_0110011;
        //mem[24] = 32'b0000000_00000_00010_100_00001_0110011;
        //mem[25] = 32'b0000000_00000_00011_100_00010_0110011;
        //mem[26] = 32'b0100000_00001_00010_000_00010_0110011;
        //mem[27] = 32'b1111101_00010_00000_001_10001_1100011; //
        //mem[28] = 32'b0000000_00100_00001_001_00001_0110011;
        //mem[29] = 32'b0000000_00001_00000_010_00000_0100011;
        //mem[30] = 32'b0000000_00000_00000_000_00000_0010011; // NOP
        //mem[31] = 32'b0000000_00010_00000_010_00000_0100011;
        //mem[32] = 32'b0000000_00000_00000_000_00000_0010011; // NOP
        //mem[33] = 32'b0000000_00001_00000_000_00000_1110011; // BREAK
    end
endmodule
